package test_pkg;

        // import the UVM package
        import uvm_pkg::*;

        // include the uvm_macros.svh
        `include "uvm_macros.svh"
        // include the tb_defs.sv
//        `include "tb_defs.sv"

        `include "ahb_xtn.sv"
        `include "ahb_agt_config.sv"
        `include "apb_agt_config.sv"
        `include "env_config.sv"
        `include "ahb_driver.sv"
        `include "ahb_monitor.sv"
        `include "ahb_sequencer.sv"
        `include "ahb_agent.sv"
        `include "ahb_agt_top.sv"
        `include "ahb_sequence.sv"

        `include "apb_xtn.sv"
        `include "apb_monitor.sv"
        `include "apb_sequencer.sv"
        `include "apb_sequence.sv"
        `include "apb_driver.sv"
        `include "apb_agent.sv"
        `include "apb_agt_top.sv"

        `include "vsequencer.sv"
        `include "vsequence.sv"
        `include "ahb2apb_sb.sv"

        `include "ahb2apb_env.sv"
        `include "ahb2apb_test.sv"
endpackage

